module pwm2(
	input enPWM, reset, clock,
	output reg PWM,
	output reg[31:0] counter
);

/* counter */
always@(posedge clock, posedge reset) begin
  //if(enPWM) begin
    if(reset)
      begin
		  counter = 0;
		  PWM = 1;
		  end 
		else 
		begin
		 if (counter >= 2)
		  PWM =0;
		  else begin
		  PWM = 1;
		  counter = counter +1; end 
		 if (counter >= 20)
		   counter = 0;
		  else
		    counter = counter +1;
		  	    
end
end


endmodule 

